module disp(input logic [3:0] count, output logic [6:0] H);
	
		always @(*)
			case(count)
				1:	H = 7'b1111001;//1
				2:	H = 7'b0100100;//2
				3:	H = 7'b0110000;//3
				4:	H = 7'b0011001;//4
				5:	H = 7'b0010010;//5
				6:	H = 7'b0000010;//6
				7:	H = 7'b1111000;//7
				8:	H = 7'b0000000;//8
				9:	H = 7'b0010000;//9
				10:H = 7'b0001000;//A
				11:H = 7'b0000011;//b
				12:H = 7'b1000110;//C
				13:H = 7'b0100001;//D
				14:H = 7'b0000110;//E
				15:H = 7'b0001110;//F
				default:H = 7'b1111111;
			endcase
endmodule